module adder(input [31:0]pc,output [31:0] newpc);
assign newpc=pc+4;
endmodule
