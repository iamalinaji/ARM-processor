module bobble(input ismet,hazard,output bobble);
assign bobble=(!ismet)||hazard;
endmodule