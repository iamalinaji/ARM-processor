module ir(input [31:0]pc,output [31:0]ir);
wire [7:0]  mem [0:65535];
    assign {mem[3], mem[2], mem[1], mem[0]}= 32'b1110_00_1_1101_0_0000_0000_000000010100; //MOV R0 ,#20 //R0 = 20
    assign{mem[7], mem[6], mem[5], mem[4]}= 32'b1110_00_1_1101_0_0000_0001_101000000001; //MOV R1 ,#4096 //R1 = 4096
     assign{mem[11],mem[10],mem[9], mem[8]}= 32'b1110_00_1_1101_0_0000_0010_000100000011; //MOV R2 ,#0xC0000000 //R2 = -1073741824
     assign{mem[15], mem[14], mem[13], mem[12]}= 32'b1110_00_0_0100_1_0010_0011_000000000010; //ADDS R3 ,R2,R2 //R3 = -2147483648 
     assign{mem[19], mem[18], mem[17], mem[16]}= 32'b1110_00_0_0101_0_0000_0100_000000000000; //ADC R4 ,R0,R0 //R4 = 41
     assign{mem[23], mem[22], mem[21], mem[20]}= 32'b1110_00_0_0010_0_0100_0101_000100000100; //SUB R5 ,R4,R4,LSL #2 //R5 = -123
     assign{mem[27], mem[26], mem[25], mem[24]}= 32'b1110_00_0_0110_0_0000_0110_000010100000; //SBC R6 ,R0,R0,LSR #1 //R6 = 10
     assign{mem[31], mem[30], mem[29], mem[28]}= 32'b1110_00_0_1100_0_0101_0111_000101000010; //ORR R7 ,R5,R2,ASR #2 //R7 = -123
     assign{mem[35], mem[34], mem[33], mem[32]}= 32'b1110_00_0_0000_0_0111_1000_000000000011; //AND R8 ,R7,R3 //R8 = -2147483648
     assign{mem[39], mem[38], mem[37], mem[36]}= 32'b1110_00_0_1111_0_0000_1001_000000000110; //MVN R9 ,R6 //R9 = -11
    assign {mem[43], mem[42], mem[41], mem[40]}= 32'b1110_00_0_0001_0_0100_1010_000000000101; //EOR R10,R4,R5 //R10 = -84
    assign {mem[47], mem[46], mem[45], mem[44]}= 32'b1110_00_0_1010_1_1000_0000_000000000110; //CMP R8 ,R6
    assign {mem[51], mem[50], mem[49], mem[48]}= 32'b0001_00_0_0100_0_0001_0001_000000000001; //ADDNE R1 ,R1,R1 //R1 = 8192
    assign {mem[55], mem[54], mem[53], mem[52]}= 32'b1110_00_0_1000_1_1001_0000_000000001000; //TST R9 ,R8
   assign {mem[59], mem[58], mem[57], mem[56]}= 32'b0000_00_0_0100_0_0010_0010_000000000010; //ADDEQ R2 ,R2,R2 //R2 = -1073741824
     assign{mem[63], mem[62], mem[61], mem[60]}= 32'b1110_00_1_1101_0_0000_0000_101100000001; //MOV R0 ,#1024 //R0 = 1024
    assign {mem[67], mem[66], mem[65], mem[64]}= 32'b1110_01_0_0100_0_0000_0001_000000000000; //STR R1 ,[R0],#0 //MEM[1024] = 8192
    assign {mem[71], mem[70], mem[69], mem[68]}= 32'b1110_01_0_0100_1_0000_1011_000000000000; //LDR R11,[R0],#0 //R11 = 8192
     assign{mem[75], mem[74], mem[73], mem[72]}= 32'b1110_01_0_0100_0_0000_0010_000000000100; //STR R2 ,[R0],#4 //MEM[1028] = -1073741824
     assign{mem[79], mem[78], mem[77], mem[76]}= 32'b1110_01_0_0100_0_0000_0011_000000001000; //STR R3 ,[R0],#8 //MEM[1032] = -2147483648
     assign{mem[83], mem[82], mem[81], mem[80]}= 32'b1110_01_0_0100_0_0000_0100_000000001101; //STR R4 ,[R0],#13 //MEM[1036] = 41
    assign {mem[87], mem[86], mem[85], mem[84]}= 32'b1110_01_0_0100_0_0000_0101_000000010000; //STR R5 ,[R0],#16 //MEM[1040] = -123
    assign {mem[91], mem[90], mem[89], mem[88]}= 32'b1110_01_0_0100_0_0000_0110_000000010100; //STR R6 ,[R0],#20 //MEM[1044] = 10
    assign {mem[95], mem[94], mem[93], mem[92]}= 32'b1110_01_0_0100_1_0000_1010_000000000100; //LDR R10,[R0],#4 //R10 = -1073741824
    assign {mem[99], mem[98], mem[97], mem[96]}= 32'b1110_01_0_0100_0_0000_0111_000000011000; //STR R7 ,[R0],#24 //MEM[1048] = -123
    assign {mem[103], mem[102], mem[101], mem[100]}= 32'b1110_00_1_1101_0_0000_0001_000000000100; //MOV R1 ,#4 //R1 = 4
    assign {mem[107], mem[106], mem[105], mem[104]}= 32'b1110_00_1_1101_0_0000_0010_000000000000; //MOV R2 ,#0 //R2 = 0
    assign {mem[111], mem[110], mem[109], mem[108]}= 32'b1110_00_1_1101_0_0000_0011_000000000000; //MOV R3 ,#0 //R3 = 0
    assign {mem[115], mem[114], mem[113], mem[112]}= 32'b1110_00_0_0100_0_0000_0100_000100000011; //ADD R4 ,R0,R3,LSL #2
    assign {mem[119], mem[118], mem[117], mem[116]}= 32'b1110_01_0_0100_1_0100_0101_000000000000; //LDR R5 ,[R4],#0
    assign {mem[123], mem[122], mem[121], mem[120]}= 32'b1110_01_0_0100_1_0100_0110_000000000100; //LDR R6 ,[R4],#4
    assign {mem[127], mem[126], mem[125], mem[124]}= 32'b1110_00_0_1010_1_0101_0000_000000000110; //CMP R5 ,R6
    assign {mem[131], mem[130], mem[129], mem[128]}= 32'b1100_01_0_0100_0_0100_0110_000000000000; //STRGT R6 ,[R4],#0
    assign {mem[135], mem[134], mem[133], mem[132]}= 32'b1100_01_0_0100_0_0100_0101_000000000100; //STRGT R5 ,[R4],#4
    assign {mem[139], mem[138], mem[137], mem[136]}= 32'b1110_00_1_0100_0_0011_0011_000000000001; //ADD R3 ,R3,#1
    assign {mem[143], mem[142], mem[141], mem[140]}= 32'b1110_00_1_1010_1_0011_0000_000000000011; //CMP R3 ,#3
    assign {mem[147], mem[146], mem[145], mem[144]}= 32'b1011_10_1_0_111111111111111111110111 ;   //BLT #-9
    assign {mem[151], mem[150], mem[149], mem[148]}= 32'b1110_00_1_0100_0_0010_0010_000000000001; //ADD R2 ,R2,
    assign {mem[155], mem[154], mem[153], mem[152]}= 32'b1110_00_0_1010_1_0010_0000_000000000001; //CMP R2 ,R1
    assign {mem[159], mem[158], mem[157], mem[156]}= 32'b1011_10_1_0_111111111111111111110011 ;   //BLT #-13
    assign {mem[163], mem[162], mem[161], mem[160]}= 32'b1110_01_0_0100_1_0000_0001_000000000000; //LDR R1 ,[R0],#0 //R1 = -2147483648
    assign {mem[167], mem[166], mem[165], mem[164]}= 32'b1110_01_0_0100_1_0000_0010_000000000100; //LDR R2 ,[R0],#4 //R2 = -1073741824
    assign {mem[171], mem[170], mem[169], mem[168]}= 32'b1110_01_0_0100_1_0000_0011_000000001000; //STR R3 ,[R0],#8 //R3 = 41
    assign {mem[175], mem[174], mem[173], mem[172]}= 32'b1110_01_0_0100_1_0000_0100_000000001100; //STR R4 ,[R0],#12 //R4 = 8192
    assign {mem[179], mem[178], mem[177], mem[176]}= 32'b1110_01_0_0100_1_0000_0101_000000010000; //STR R5 ,[R0],#16 //R5 = -123
    assign {mem[183], mem[182], mem[181], mem[180]}= 32'b1110_01_0_0100_1_0000_0110_000000010100; //STR R6 ,[R0],#20 //R4 = 10
    assign {mem[187], mem[186], mem[185], mem[184]}= 32'b1110_10_1_0_111111111111111111111111 ;   //B #-1
assign ir={mem[pc+3],mem[pc+2],mem[pc+1],mem[pc]};
endmodule